module key_module128(
input [255:0] key,
input [1:0] Algorithm,
input [3:0] i,
output reg [127:0] out
);

wire [255:0] keyin1;
wire [255:0] keyin2;
wire [255:0] keyin3;
wire [255:0] keyin4;
wire [255:0] keyin5;
wire [255:0] keyin6;
wire [255:0] keyin7;
wire [255:0] keyin8;
wire [255:0] keyin9;
wire [255:0] keyin10;

wire [1408:0] array; 
wire [255:0]key_exp_out1;
wire [255:0]key_exp_out2;
wire [255:0]key_exp_out3;
wire [255:0]key_exp_out4;
wire [255:0]key_exp_out5;
wire [255:0]key_exp_out6;
wire [255:0]key_exp_out7;
wire [255:0]key_exp_out8;
wire [255:0]key_exp_out9;
wire [255:0]key_exp_out10;

//0 original 1128 key
assign array[1408:1280]=key[255:128];
//1
assign keyin1=key;
Key_Expansion_new  singleKeyExpansionInst1 (keyin1,4'h1,2'b00,key_exp_out1);
assign array[1279:1152]=key_exp_out1[255:128];
//2
assign keyin2=key_exp_out1;
Key_Expansion_new  singleKeyExpansionInst2 (keyin2,4'h2,2'b00,key_exp_out2);
assign array[1151:1024]=key_exp_out2[255:128];
//3
assign keyin3=key_exp_out2;
Key_Expansion_new  singleKeyExpansionInst3 (keyin3,4'h3,2'b00,key_exp_out3);
assign array[1023:896]=key_exp_out3[255:128];
//4
assign keyin4=key_exp_out3;
Key_Expansion_new  singleKeyExpansionInst4 (keyin4,4'h4,2'b00,key_exp_out4);
assign array[895:768]=key_exp_out4[255:128];
//5
assign keyin5=key_exp_out4;
Key_Expansion_new  singleKeyExpansionInst5 (keyin5,4'h5,2'b00,key_exp_out5);
assign array[767:640]=key_exp_out5[255:128];
//6
assign keyin6=key_exp_out5;
Key_Expansion_new  singleKeyExpansionInst6 (keyin6,4'h6,2'b00,key_exp_out6);
assign array[639:512]=key_exp_out6[255:128];
//7
assign keyin7=key_exp_out6;
Key_Expansion_new  singleKeyExpansionInst7 (keyin7,4'h7,2'b00,key_exp_out7);
assign array[511:384]=key_exp_out7[255:128];
//8
assign keyin8=key_exp_out7;
Key_Expansion_new  singleKeyExpansionInst8 (keyin8,4'h8,2'b00,key_exp_out8);
assign array[383:256]=key_exp_out8[255:128];
//9
assign keyin9=key_exp_out8;
Key_Expansion_new  singleKeyExpansionInst9 (keyin9,4'h9,2'b00,key_exp_out9);
assign array[255:128]=key_exp_out9[255:128];
//10
assign keyin10=key_exp_out9;
Key_Expansion_new  singleKeyExpansionInst10 (keyin10,4'ha,2'b00,key_exp_out10);
assign array[127:0]=key_exp_out10[255:128];

always@(*)begin
//originla key
if(i==0)begin
out=array[1408:1280];
end
if(i==1)begin
out=array[1280:1152];
end
if(i==2)begin
out=array[1151:1024];
end
if(i==3)begin
out=array[1023:896];
end
if(i==4)begin
out=array[895:768];
end
if(i==5)begin
out=array[767:640];
end
if(i==6)begin
out=array[639:512];
end
if(i==7)begin
out=array[511:384];
end
if(i==8)begin
out=array[383:256];
end
if(i==9)begin
out=array[255:128];
end
if(i==10)begin
out=array[127:0];
end
end

endmodule
